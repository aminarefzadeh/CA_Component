module datapath(input pop,push,memorywrite,memoryread,writeReg,selRR2,selALU2,selpc,ldz,ldc,selz,selc,input [1:0] selWD,selRet,input  [2:0]ALUfn,input clk,rst, output reg ze,c,output reg[5:0] code);
  wire [11:0] pc_1 , ret;
  stack Stack(pc_1,push,pop,clk,rst,ret);
  wire[11:0] f_pc,next_pc;
  wire [18:0] ins;
  mux3_12 pc_ret(f_pc , ret , ins[11:0] , selRet ,next_pc);
  wire[11:0] pc;
  pc PC(next_pc ,clk,rst,pc);
  instructionMem IM(pc,rst,ins);
  wire [11:0]extended;
  signExtender Ex(ins[7:0], extended );
  adder_1 In(pc ,pc_1);
  wire[11:0] apc;
  adder Add(pc_1 , extended , apc);
  mux2_12 pc1_apc(pc_1 , apc , selpc , f_pc);
  wire [2:0] RR2;
  mux2_3 sel_RR2(ins[7:5] , ins[13:11] , selRR2, RR2);
  wire [7:0] Out,RD,ALUOut,WD;
  mux3 sel_WD( ALUOut,RD,Out, selWD,WD);
  wire[7:0] RD1,RD2;
  registerFile RF(ins[10:8],RR2,ins[13:11],WD,writeReg,clk,rst,RD1,RD2);
  wire[7:0] ALU2;
  mux2_8 sel_ALU2(ins[7:0] , RD2, selALU2,ALU2);
  wire zero,carry;
  alu Alu(ALUfn ,RD1,ALU2 ,c ,ALUOut ,zero,carry);
  wire shc,shz;
  shiftReg Shr(RD1,ins[7:5],ins[15:14],Out,shc,shz);
  wire ff1;
  mux2_1 sel_z(zero,shz,selz , ff1);
  ff ff_z(ff1,ldz,clk,rst,ze);
  wire ff2;
  mux2_1 sel_c(carry,shc,selc , ff2);
  ff ff_c(ff2,ldc,clk,rst,c);
  memory Mem(ALUOut,RD2,clk,memorywrite,memoryread,RD);
  assign code = ins[18:13];
endmodule